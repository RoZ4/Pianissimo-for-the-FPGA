`define STARTSCREEN 5'd0
`define RECORD 5'd1
`define PLAYBACK 5'd2
`define RESTARTPLAYBACK 5'd3
`define NUMBEROFKEYBOARDINPUTS 30