/* This module implements the VGA controller. It assumes a 25MHz clock is supplied as input.
 * General approach:
 * Go through each line of the screen and read the colour each pixel on that line should have from
 * the Video memory. To do that for each (x,y) pixel on the screen convert (x,y) coordinate to
 * a memory_address at which the pixel colour is stored in Video memory. Once the pixel colour is
 * read from video memory its brightness is first increased before it is forwarded to the VGA DAC.
 */
module vga_controller(vga_clock, resetn, pixel_colour, memory_address, 
		VGA_R, VGA_G, VGA_B,
		VGA_HS, VGA_VS, VGA_BLANK_N,
		VGA_SYNC_N, VGA_CLK);
	
	/* Colour depth and screen resolution parameters; see the vga_adapter module for descriptions
    * of each parameter. */
	parameter BITS_PER_COLOUR_CHANNEL = 1;
	parameter MONOCHROME = "FALSE";
	parameter RESOLUTION = "320x240";
	//--- Timing parameters.
	/* Recall that the VGA specification requires a few more rows and columns are drawn
	 * when refreshing the screen than are actually present on the screen. This is necessary to
	 * generate the vertical and the horizontal syncronization signals. If you wish to use a
	 * display mode other than 640x480 you will need to modify the parameters below as well
	 * as change the frequency of the clock driving the monitor (VGA_CLK).
	 */
	parameter C_VERT_NUM_PIXELS  = 11'd480;
	parameter C_VERT_SYNC_START  = 11'd493;
	parameter C_VERT_SYNC_END    = 11'd494; //(C_VERT_SYNC_START + 2 - 1); 
	parameter C_VERT_TOTAL_COUNT = 11'd525;

	parameter C_HORZ_NUM_PIXELS  = 11'd640;
	parameter C_HORZ_SYNC_START  = 11'd659;
	parameter C_HORZ_SYNC_END    = 11'd754; //(C_HORZ_SYNC_START + 96 - 1); 
	parameter C_HORZ_TOTAL_COUNT = 11'd800;	
		
	/*****************************************************************************/
	/* Declare inputs and outputs.                                               */
	/*****************************************************************************/
	
	input vga_clock, resetn;
	input [((MONOCHROME == "TRUE") ? (0) : (BITS_PER_COLOUR_CHANNEL*3-1)):0] pixel_colour;
	output [((RESOLUTION == "320x240") ? (16) : (14)):0] memory_address;
	output reg [7:0] VGA_R;
	output reg [7:0] VGA_G;
	output reg [7:0] VGA_B;
	output reg VGA_HS;
	output reg VGA_VS;
	output reg VGA_BLANK_N;
	output VGA_SYNC_N, VGA_CLK;
	
	/*****************************************************************************/
	/* Local Signals.                                                            */
	/*****************************************************************************/
	
	reg VGA_HS1;
	reg VGA_VS1;
	reg VGA_BLANK1; 
	reg [9:0] xCounter, yCounter;
	wire xCounter_clear;
	wire yCounter_clear;
	wire vcc;
	
	reg [((RESOLUTION == "320x240") ? (8) : (7)):0] x; 
	reg [((RESOLUTION == "320x240") ? (7) : (6)):0] y;	
	/* Inputs to the converter. */
	
	/*****************************************************************************/
	/* Controller implementation.                                                */
	/*****************************************************************************/

	assign vcc =1'b1;
	
	/* A counter to scan through a horizontal line. */
	always @(posedge vga_clock or negedge resetn)
	begin
		if (!resetn)
			xCounter <= 10'd0;
		else if (xCounter_clear)
			xCounter <= 10'd0;
		else
		begin
			xCounter <= xCounter + 1'b1;
		end
	end
	assign xCounter_clear = (xCounter == (C_HORZ_TOTAL_COUNT-1));

	/* A counter to scan vertically, indicating the row currently being drawn. */
	always @(posedge vga_clock or negedge resetn)
	begin
		if (!resetn)
			yCounter <= 10'd0;
		else if (xCounter_clear && yCounter_clear)
			yCounter <= 10'd0;
		else if (xCounter_clear)		//Increment when x counter resets
			yCounter <= yCounter + 1'b1;
	end
	assign yCounter_clear = (yCounter == (C_VERT_TOTAL_COUNT-1)); 
	
	/* Convert the xCounter/yCounter location from screen pixels (640x480) to our
	 * local dots (320x240 or 160x120). Here we effectively divide x/y coordinate by 2 or 4,
	 * depending on the resolution. */
	always @(*)
	begin
		if (RESOLUTION == "320x240")
		begin
			x = xCounter[9:1];
			y = yCounter[8:1];
		end
		else
		begin
			x = xCounter[9:2];
			y = yCounter[8:2];
		end
	end
	
	/* Change the (x,y) coordinate into a memory address. */
	vga_address_translator controller_translator(
					.x(x), .y(y), .mem_address(memory_address) );
		defparam controller_translator.RESOLUTION = RESOLUTION;


	/* Generate the vertical and horizontal synchronization pulses. */
	always @(posedge vga_clock)
	begin
		//- Sync Generator (ACTIVE LOW)
		VGA_HS1 <= ~((xCounter >= C_HORZ_SYNC_START) && (xCounter <= C_HORZ_SYNC_END));
		VGA_VS1 <= ~((yCounter >= C_VERT_SYNC_START) && (yCounter <= C_VERT_SYNC_END));
		
		//- Current X and Y is valid pixel range
		VGA_BLANK1 <= ((xCounter < C_HORZ_NUM_PIXELS) && (yCounter < C_VERT_NUM_PIXELS));	
	
		//- Add 1 cycle delay
		VGA_HS <= VGA_HS1;
		VGA_VS <= VGA_VS1;
		VGA_BLANK_N <= VGA_BLANK1;	
	end
	
	/* VGA sync should be 1 at all times. */
	assign VGA_SYNC_N = vcc;
	
	/* Generate the VGA clock signal. */
	assign VGA_CLK = vga_clock;
	
	/* Brighten the colour output. */
	// The colour input is first processed to brighten the image a little. Setting the top
	// bits to correspond to the R,G,B colour makes the image a bit dull. To brighten the image,
	// each bit of the colour is replicated through the 10 DAC colour input bits. For example,
	// when BITS_PER_COLOUR_CHANNEL is 2 and the red component is set to 2'b10, then the
	// VGA_R input to the DAC will be set to 10'b1010101010.
	
	integer index;
	integer sub_index;
	
	wire on_screen;
	
	assign on_screen = (({1'b0, xCounter} >= 0) & ({1'b0, xCounter} < C_HORZ_NUM_PIXELS+2) & ({1'b0, yCounter} < C_VERT_NUM_PIXELS));
	
	always @(pixel_colour or on_screen)
	// Translate 3bit colour to custom palette (3 shades of blue, 3 shades of red, black, white 256/3 = 85.333)
	begin
		VGA_R <= 'b0;
		VGA_G <= 'b0;
		VGA_B <= 'b0;
		if (MONOCHROME == "FALSE") begin
			case(pixel_colour)
				'd0: begin 				  // WHITE
					VGA_R <= 8'b11111111;
					VGA_G <= 8'b11111111;
					VGA_B <= 8'b11111111;
					
					end
				'd1: begin 				  // BLUE
					VGA_R <= 8'b00000000;
					VGA_G <= 8'b00000000;
					VGA_B <= 8'b11111111;
					end
				'd2: begin
					VGA_R <= 8'b11010101; //213
					VGA_G <= 8'b11010101;
					VGA_B <= 8'b11111111;
					end
				'd3: begin
					VGA_R <= 8'b10101010; //170
					VGA_G <= 8'b10101010;
					VGA_B <= 8'b11111111;
					end
				'd4: begin 				  
					VGA_R <= 8'b01111111; // 127
					VGA_G <= 8'b11111111;
					VGA_B <= 8'b11111111;
					end
				'd5: begin
					VGA_R <= 8'b01010100; // 84
					VGA_G <= 8'b01010100;
					VGA_B <= 8'b11111111;
					end
				'd6: begin
					VGA_R <= 8'b00101011; //43
					VGA_G <= 8'b00101011;
					VGA_B <= 8'b11111111;
					end
				'd7: begin 				  // BLACK
					VGA_R <= 8'b00000000;
					VGA_G <= 8'b00000000;
					VGA_B <= 8'b00000000;
					end
				// 'd0: begin 				  // BLACK
				// 	VGA_R <= 8'b00000000;
				// 	VGA_G <= 8'b00000000;
				// 	VGA_B <= 8'b00000000;
				// 	end
				// 'd1: begin 				  // BLUE
				// 	VGA_R <= 8'b00000000;
				// 	VGA_G <= 8'b00000000;
				// 	VGA_B <= 8'b11111111;
				// 	end
				// 'd2: begin
				// 	VGA_R <= 8'b10101100; //172
				// 	VGA_G <= 8'b10101100;
				// 	VGA_B <= 8'b11111111;
				// 	end
				// 'd3: begin
				// 	VGA_R <= 8'b01010110; //86
				// 	VGA_G <= 8'b01010110;
				// 	VGA_B <= 8'b11111111;
				// 	end
				// 'd4: begin 				  // RED
				// 	VGA_R <= 8'b11111111;
				// 	VGA_G <= 8'b00000000;
				// 	VGA_B <= 8'b00000000;
				// 	end
				// 'd5: begin
				// 	VGA_R <= 8'b11111111;
				// 	VGA_G <= 8'b10101100;
				// 	VGA_B <= 8'b10101100;
				// 	end
				// 'd6: begin
				// 	VGA_R <= 8'b11111111;
				// 	VGA_G <= 8'b01010110;
				// 	VGA_B <= 8'b01010110;
				// 	end
				// 'd7: begin 				  // WHITE
				// 	VGA_R <= 8'b11111111;
				// 	VGA_G <= 8'b11111111;
				// 	VGA_B <= 8'b11111111;
				// 	end
			endcase
		end
	end

			

	/*
	begin		
		VGA_R <= 'b0;
		VGA_G <= 'b0;
		VGA_B <= 'b0;
		if (MONOCHROME == "FALSE")
		begin
			for (index = 8-BITS_PER_COLOUR_CHANNEL; index >= 0; index = index - BITS_PER_COLOUR_CHANNEL)
			begin
				for (sub_index = BITS_PER_COLOUR_CHANNEL - 1; sub_index >= 0; sub_index = sub_index - 1)
				begin
					VGA_R[sub_index+index] <= on_screen & pixel_colour[sub_index + BITS_PER_COLOUR_CHANNEL*2];
					VGA_G[sub_index+index] <= on_screen & pixel_colour[sub_index + BITS_PER_COLOUR_CHANNEL];
					VGA_B[sub_index+index] <= on_screen & pixel_colour[sub_index];
				end
			end	
		end
		else
		begin
			for (index = 0; index < 8; index = index + 1)
			begin
				VGA_R[index] <= on_screen & pixel_colour[0:0];
				VGA_G[index] <= on_screen & pixel_colour[0:0];
				VGA_B[index] <= on_screen & pixel_colour[0:0];
			end	
		end
	end
	*/

endmodule
